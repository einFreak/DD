library IEEE; 
use IEEE.STD_LOGIC_1164.all;
entity module is
  port(clk, reset, a, b: in  STD_LOGIC;
    q: out STD_LOGIC);
end;

architecture arch of module is
--##INSERT YOUR CODE HERE 
  --type statetype is (S0, S1, S2);
  --signal state, nstate: statetype;
begin
  
  
--##INSERT YOUR CODE HERE END
end;
