library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity MODULE is
  port( CLK, RESET: in std_logic;
        segments: out std_logic_vector(6 downto 0)
      );
end MODULE;

architecture arch of MODULE is
--##INSERT YOUR CODE HERE
 
--##INSERT YOUR CODE HERE END

end;
