library ieee; 
use ieee.std_logic_1164.all; 
--use ieee.numeric_std.all;     
use ieee.std_logic_unsigned.all;   

entity module is 
  port( CLK, RESET: in std_logic; 
    MODE: in  std_logic_vector(1 downto 0); 
    Q: out std_logic_vector(3 downto 0)); 
end; 
 
architecture arch of module is 
--##INSERT YOUR CODE HERE 
  --signal Q_INT : std_logic_vector(3 downto 0); --local signal 
begin 

--##INSERT YOUR CODE HERE 
end; 
